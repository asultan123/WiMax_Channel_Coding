library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity wimax_tb is   
end  wimax_tb;
architecture behav of wimax_tb is
component wimax is
   port(
      clk_m, clk2_m, reset_m: in std_logic;
	  ready_m : in std_logic;
	  data_in_m : in std_logic;
	  seed_m : in std_logic_vector(0 to 14);
	  valid_m: out std_logic;
	  data_out0_m, data_out1_m: out std_logic_vector(15 downto 0)
   );
end component ;

signal  clk1:  std_logic := '0';
signal clk2: std_logic := '1';
signal  reset:  std_logic;
signal  ready, data_in:  std_logic;
signal seed :  std_logic_vector(0 to 14);
signal valid:  std_logic;
signal data_out0: std_logic_vector (15 downto 0);
signal data_out1: std_logic_vector (15 downto 0);
signal input: std_logic_vector(0 to 95) := x"ACBCD2114DAE1577C6DBF4C9";
------
signal rightI:std_logic_vector(959 downto 0):="011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001";
signal rightQ:std_logic_vector(959 downto 0):="110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100";
signal zerosI,zerosQ:std_logic_vector(959 downto 0);


constant PERIOD2: time := 10 ns;
constant PERIOD1: time := 20 ns;
begin

uut: wimax 
	port map(
    clk_m	=> clk1,
	clk2_m => clk2,
    reset_m	=> reset,
    ready_m	=> ready,
	seed_m => seed,
    data_in_m	 => data_in,
    valid_m => valid,
    data_out0_m => data_out0,
	data_out1_m => data_out1
    );
	

 clk1 <= not clk1 after PERIOD1/2;
 clk2 <= not clk2 after PERIOD2/2;

 
 stimulus : process 
 
	begin
	reset <= '1';
	wait for (PERIOD1); reset <='0';
	wait for (PERIOD1);
	ready <= '1';
	seed <= "011011100010101";
	for i in 0 to 959 loop
		data_in <= input(i mod 96);
		wait for (1*PERIOD1);
    end loop;
	ready <= '0';
	wait;
	
	

end  process stimulus;



process
variable error_status:boolean; 
begin
wait until (valid = '1');
for z in 959 downto 0 loop
		
		wait for (PERIOD2);
  
	 
		if (data_out0="0101101001111111") then
		zerosI(z)<='1'; 
		else 
		zerosI(z)<='0';
		end if;
		if (data_out1="0101101001111111") then
		zerosQ(z)<='1'; 
		else 
		zerosQ(z)<='0';
		end if;
		wait for(PERIOD2);
		
	
end loop;


if((zerosI=rightI) and (zerosQ=rightQ)) then 
	error_status := true;
else
	error_status := false;
end if;
assert error_status
report "test failed."
severity note;
	
end process;

end behav;             
                                       