library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity modulator_tb is
end modulator_tb;

architecture modulator_tb_arch of modulator_tb is 
component modulator
port(
	reset, clk, en:in std_logic;
	d:in std_logic;
	valid:out std_logic;
	I:out std_logic_vector(15 downto 0);
	Q:out std_logic_vector(15 downto 0)
	);
end component;

signal clk:std_logic:='1';
signal reset, en, d, valid:std_logic:='0';
signal I, Q:std_logic_vector(15 downto 0);
signal input_test:std_logic_vector(191 downto 0):=x"4B047DFA42F2A5D5F61C021A5851E9A309A24FD58086BD1E";												
signal rightI:std_logic_vector(959 downto 0):="011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001011011010000001101110011110000000001100111111011001100100110111011101111010000001111110110001001";
signal rightQ:std_logic_vector(959 downto 0):="110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100110011111001000011100010001101110010110111101100110111110001001011010010110001110111011000011100";
signal zerosI,zerosQ:std_logic_vector(959 downto 0);
signal flag:std_logic := '0';
constant PERIOD:time:=10 ns;

begin
dut:modulator port map(reset=>reset, clk=>clk, en=>en, d=>d, valid=>valid, I=>I, Q=>Q);

clk<=not clk after PERIOD/2;

stimulus:process
variable error_status:boolean;

variable mimi: integer:=1919;
begin
reset  <= '1'; wait for 0.7*PERIOD; 
reset  <= '0'; 
en<='1'; 

for z in 959 downto 0 loop
  d<=input_test(mimi mod 192);

	wait for PERIOD;
	flag <= '0';
	mimi := mimi-1;
	
	
d<=input_test(mimi mod 192);	

	wait for PERIOD;
	flag <= not (flag);
	mimi:= mimi-1;
	
end loop;

en<='0'; wait for 2*PERIOD;


if((zerosI=rightI) and (zerosQ=rightQ)) then 
	error_status := true;
else
	error_status := false;
end if;
assert error_status
report "test failed."
severity failure;
wait;
end process stimulus;

process 

variable  k:integer:=959;

begin
wait on flag;
if (flag = '1') then 
	if (I="0101101001111111") then
	zerosI(k)<='1'; 
	else 
	zerosI(k)<='0';
	end if;
	if (Q="0101101001111111") then
	zerosQ(k)<='1'; 
	else 
	zerosQ(k)<='0';
	end if;
	
k := k - 1;

end if;

end process;

end modulator_tb_arch;
